--/////////////////////////////////////////////////////////////////////////////////////////
-- Company: Digilent Inc.
-- Engineer: Josh Sackos
-- 
-- Create Date:    07/26/2012
-- Module Name:    PmodACL_Demo
-- Project Name: 	 PmodACL_Demo
-- Target Devices: Nexys3
-- Tool versions:  ISE 14.1
-- Description: This is a demo for the Digilent PmodACL.  The SW inputs are
--					 used to select either the x-axis, y-axis, or z-axis data for
--					 display, and RST is used to reset the demo.
--
--					 There are four main components in this module, SPIcomponent, sel_Data,
--					 ClkDiv_5Hz, and ssdCtrl.  A START signal is generated by the ClkDiv_5Hz
--					 component, this signal is used to initiate a data transfer between the
--					 PmodACL and the Nexys3.
--
--					 SPIcomponent receives the START signal, configures the PmodACL, and then
--					 receives data pertaining to all three axes.  The data is made available
--					 to the rest of the design on the xAxis, yAxis, and zAxis outputs.
--
--					 These outputs are then sent into the sel_Data component with the the status
--					 of switches SW1 and SW0 on the Nexys3. Depending on the configuration of
--					 these switches, one of the axes data will be selected for display on the
--					 seven segment display. The selected data is converted from 2's compliment
--					 to magnitude, and is then sent to the ssdCtrl where it is converted to a "g"
--					 value and displayed on the SSD with hundredths precision.
--
--					 To select an axis for display configure SW1 and SW0 on the Nexys3 as
--					 shown below.  LED LD0 will illuminate when the x-axis is selected,
--					 LD1 for y-aixs, and LD2 for z-axis.
--
--							SW1	SW0	|	SSD Output	|	LD2	|	LD1	|	LD0
--							------------------------------------------------------
--							off	off	|	x-axis		|	off	|	off	|	on
--							off	on		|	y-axis		|	off	|	on		|	off
--							on		on		|	x-axis		|	off	|	off	|	on
--							on		off	|	z-axis		|	on		|	off	|	off
--

--  Inputs:
--		CLK				Onboard system clock
--		RST				Resets the demo
--		SW<0>				Selects y-axis data for display
--		SW<1>				Selects z-axis data for display
--		SDI				Serial Data In
--
--  Outputs:
--		SDO				Serial Data Out
--		SCLK				Serial Clock
--		SS					Slave Select
--		AN					Anodes on SSD
--		SEG				Cathodes on SSD
--		DOT				Cathode for decimal on SSD
--		LED				LEDs on Nexys3
--
-- Revision History: 
-- 						Revision 0.01 - File Created (Josh Sackos)
--/////////////////////////////////////////////////////////////////////////////////////////
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_arith.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- ====================================================================================
-- 										  Define Module
-- ====================================================================================
entity PmodACL_Demo is
    Port ( CLK : in  STD_LOGIC;
           RST : in  STD_LOGIC;
           SW : in  STD_LOGIC_VECTOR (2 downto 0);
           SDI : in  STD_LOGIC;
           SDO : out  STD_LOGIC;
           SCLK : out  STD_LOGIC;
           SS : out  STD_LOGIC;
           AN : out  STD_LOGIC_VECTOR (3 downto 0);
           SEG : out  STD_LOGIC_VECTOR (6 downto 0);
           DOT : out  STD_LOGIC;
           LED : out  STD_LOGIC_VECTOR (2 downto 0);
			  
			  LV : in  STD_LOGIC_VECTOR (1 downto 0);
			  
			  --vga outputs
			  rgb_out:  out std_logic_vector(7 downto 0);
			  hs_out: out std_logic;
			  vs_out: out std_logic;
			  
			  --for debugging
			  Data: out STD_LOGIC_VECTOR (7 downto 0);
			  
			  s_x : out STD_LOGIC_VECTOR (1 downto 0);
			  s_y : out STD_LOGIC_VECTOR (1 downto 0);
			  --s_l : out STD_LOGIC_VECTOR (1 downto 0);
			  --s_r : out STD_LOGIC_VECTOR (1 downto 0);
			  
			  x_dir : out STD_LOGIC;
			  y_dir : out STD_LOGIC
	);
end PmodACL_Demo;

architecture Behavioral of PmodACL_Demo is


--  ===================================================================================
-- 							  				  Components
--  ===================================================================================

		-- **********************************************
		-- 		 			 Select Data
		-- **********************************************
		component sel_Data Port(
					CLK : in  STD_LOGIC;
					RST : in  STD_LOGIC;
					SW : in STD_LOGIC_VECTOR(1 downto 0);
					xAxis : in  STD_LOGIC_VECTOR (9 downto 0);
					yAxis : in  STD_LOGIC_VECTOR (9 downto 0);
					zAxis : in  STD_LOGIC_VECTOR (9 downto 0);
					DOUT : out  STD_LOGIC_VECTOR (9 downto 0);
					LED : out  STD_LOGIC_VECTOR (2 downto 0)
		);
		end component;

		-- **********************************************
		-- 		 Seven Segment Display Controller
		-- **********************************************
		component SPIcomponent
			Port ( CLK : in  STD_LOGIC;
					 RST : in  STD_LOGIC;
					 START : in STD_LOGIC;
					 SDI : in  STD_LOGIC;
					 SDO : out  STD_LOGIC;
					 SCLK : out  STD_LOGIC;
					 SS : out  STD_LOGIC;
					 xAxis : out STD_LOGIC_VECTOR(9 downto 0);
					 yAxis : out STD_LOGIC_VECTOR(9 downto 0);
					 zAxis : out STD_LOGIC_VECTOR(9 downto 0)
			 );
		end component;

		-- **********************************************
		-- 		 Seven Segment Display Controller
		-- **********************************************
--		component ssdCtrl
--			 Port ( CLK : in  STD_LOGIC;
--					  RST : in  STD_LOGIC;
--					  DIN : in  STD_LOGIC_VECTOR (9 downto 0);
--					  AN : out  STD_LOGIC_VECTOR (3 downto 0);
--					  SEG : out  STD_LOGIC_VECTOR (6 downto 0);
--					  DOT : out STD_LOGIC
--			 );
--		end component;

		-- **********************************************
		-- 				5Hz Clock Divider
		-- **********************************************
		component ClkDiv_5Hz
			Port (  CLK : in  STD_LOGIC;
					  RST : in STD_LOGIC;
					  CLKOUT : inout STD_LOGIC);
		end component;
		
		-- **********************************************
		-- 				Speed Calculator Module
		-- **********************************************
		component speedCalculator
			Port (  --xAxis :  in  STD_LOGIC_VECTOR (9 downto 0);
					  --yAxis :  in  STD_LOGIC_VECTOR (9 downto 0);
					  xAxis :  in  STD_LOGIC_VECTOR (9 downto 0);
					  yAxis :  in  STD_LOGIC_VECTOR (9 downto 0);
					  sp_x : out STD_LOGIC_VECTOR(1 downto 0);
					  sp_y : out STD_LOGIC_VECTOR(1 downto 0)
			);
		end component;
		
		component VGAOutput
			Port (  
						v_dir : in STD_LOGIC;
						h_dir : in STD_LOGIC;
						sp_v : in STD_LOGIC_VECTOR(1 downto 0);
						sp_h : in STD_LOGIC_VECTOR(1 downto 0);
						
						clk100_in: in std_logic;
						rst : in std_logic;
						lv : in STD_LOGIC_VECTOR(1 downto 0);

						rgb_out:  out std_logic_vector(7 downto 0);
						hs_out: out std_logic;
						vs_out: out std_logic
			);
		end component;



-- ====================================================================================
-- 							       Signals and Constants
-- ====================================================================================

		signal xAxis : STD_LOGIC_VECTOR(9 downto 0);		-- x-axis data from PmodACL
		signal yAxis : STD_LOGIC_VECTOR(9 downto 0);		-- y-axis data from PmodACL
		signal zAxis : STD_LOGIC_VECTOR(9 downto 0);		-- z-axis data from PmodACL

		signal selData : STD_LOGIC_VECTOR(9 downto 0);	-- Data selected to display

		signal START : STD_LOGIC;								-- Data Transfer Request Signal

		signal spd_x : STD_LOGIC_VECTOR(1 downto 0) := "00";
		signal spd_y : STD_LOGIC_VECTOR(1 downto 0) := "00";
		--signal spd_l : STD_LOGIC_VECTOR(1 downto 0) := "00";
		--signal spd_r : STD_LOGIC_VECTOR(1 downto 0) := "00";
		
--  ===================================================================================
-- 							  				Implementation
--  ===================================================================================
begin

			-------------------------------------------------
			--	Select Display Data and Convert to Magnitude
			-------------------------------------------------
			SDATA : sel_Data port map(
							CLK=>CLK,
							RST=>RST,
							SW=>SW(1 downto 0),
							xAxis=>xAxis,
							yAxis=>yAxis,
							zAxis=>zAxis,
							DOUT=>selData,
							LED=>LED
			);

			-------------------------------------------------
			--		 			 Interfaces PmodACL
			-------------------------------------------------
			SPI : SPIcomponent port map(
							CLK=>CLK,
							RST=>RST,
							START=>START,
							SDI=>SDI,
							SDO=>SDO,
							SCLK=>SCLK,
							SS=>SS,
							xAxis=>xAxis,
							yAxis=>yAxis,
							zAxis=>zAxis
			);

			-------------------------------------------------
			--		 	 Formats Data and Displays on SSD
			-------------------------------------------------
--			Disp : ssdCtrl port map(
--							CLK=>CLK,
--							RST=>RST,
--							DIN=>selData(9 downto 0),
--							AN=>AN,
--							SEG=>SEG,
--							DOT=>DOT
--			);

			-------------------------------------------------
			--	 Generates a 5Hz Data Transfer Request Signal
			-------------------------------------------------
			genStart : ClkDiv_5Hz port map(
							CLK=>CLK,
							RST=>RST,
							CLKOUT=>START
			);
			
			calcSpeeds : speedCalculator port map (
							xAxis=>xAxis(9 downto 0),
							yAxis=>yAxis(9 downto 0),
							sp_x=>spd_x,
							sp_y=>spd_y
							--sp_l=>spd_l,
							--sp_r=>spd_r
			);
			
			printScreen: VGAOutput port map (
							v_dir=>xAxis(9),
							h_dir=>yAxis(9),
							sp_v=>spd_x(1 downto 0),
							sp_h=>spd_y(1 downto 0),
							
							clk100_in=>CLK,
							rst=>RST,
							lv => LV,
							
							rgb_out=>rgb_out,
							hs_out=>hs_out,
							vs_out=>vs_out
			);
			
			process 
			begin
			
--			if SW(2) = '1' then
--				Data(7) <= xAxis(9);
--				Data(6 downto 5) <= spd_x(1 downto 0);
--				Data(4 downto 3) <= "00";
--				Data(2) <= yAxis(9);
--				Data(1 downto 0) <= spd_y(1 downto 0);
--			else 
--				if SW(1 downto 0) = "00" then
--					Data <= xAxis(7 downto 0);
--				elsif SW(1 downto 0) = "01" then 
--					Data <= yAxis(7 downto 0);
--				else
--					Data <= selData(7 downto 0);
--				end if;
--			end if;
			
--			-- old debug
--			--s_u <= "00";
--			s_x <= spd_x(1 downto 0);
--			--s_l <= "00";
--			s_y <= spd_y(1 downto 0);
--			
--			x_dir <= xAxis(9);
--			y_dir <= yAxis(9);
--			
			end process;
end Behavioral;

